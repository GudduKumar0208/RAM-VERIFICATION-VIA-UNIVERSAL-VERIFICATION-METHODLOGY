class ram_config extends uvm_object;

`uvm_object_utils(ram_config)

function new(string name="ram_config");
super.new(name);

endfunction

bit scoreboard=0;

endclass